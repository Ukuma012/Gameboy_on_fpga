// top module

module UGB(
    input logic pin_clk,
    input logic pin_n_reset
);